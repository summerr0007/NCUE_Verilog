module sort8_pipe_2(clk,rst,x0,x1,x2,x3,x4,x5,x6,x7,y0,y1,y2,y3,y4,y5,y6,y7);
	input clk, rst;
	input [7:0] x0,x1,x2,x3,x4,x5,x6,x7;
	output [7:0] y0,y1,y2,y3,y4,y5,y6,y7;
	wire [7:0] a0,b0,c0,d0,e0,f0;
	wire [7:0] a1,b1,c1,d1,e1,f1;
	wire [7:0] a2,b2,c2,d2,e2,f2;
	wire [7:0] a3,b3,c3,d3,e3,f3;
	wire [7:0] a4,b4,c4,d4,e4,f4;
	wire [7:0] a5,b5,c5,d5,e5,f5;
	wire [7:0] a6,b6,c6,d6,e6,f6;
	wire [7:0] a7,b7,c7,d7,e7,f7;
	dff r00 (x0,clk,rst,a0);
	dff r01 (x1,clk,rst,a1);
	dff r02 (x2,clk,rst,a2);
	dff r03 (x3,clk,rst,a3);
	dff r04 (x4,clk,rst,a4);
	dff r05 (x5,clk,rst,a5);
	dff r06 (x6,clk,rst,a6);
	dff r07 (x7,clk,rst,a7);
	sort4_pipe inst0(clk,rst,a0,a1,a2,a3,b0,b1,b2,b3);
	sort4_pipe inst1(clk,rst,a4,a5,a6,a7,b4,b5,b6,b7);
	dff r10 (b0,clk,rst,c0);
	dff r11 (b1,clk,rst,c1);
	dff r12 (b2,clk,rst,c2);
	dff r13 (b3,clk,rst,c3);
	dff r14 (b4,clk,rst,c4);
	dff r15 (b5,clk,rst,c5);
	dff r16 (b6,clk,rst,c6);
	dff r17 (b7,clk,rst,c7);
	sort4_pipe inst2(clk,rst,c0,c1,c4,c5,d0,d1,d8,d9);
	sort4_pipe inst3(clk,rst,c2,c3,c6,c7,d10,d11,d6,d7);
	dff r20 (d0,clk,rst,e0);
	dff r21 (d1,clk,rst,e1);
	dff r22 (d8,clk,rst,e8);
	dff r23 (d9,clk,rst,e9);
	dff r24 (d10,clk,rst,e10);
	dff r25 (d11,clk,rst,e11);
	dff r26 (d6,clk,rst,e6);
	dff r27 (d7,clk,rst,e7);
	sort4_pipe inst4(clk,rst,e8,e9,e10,e11,f2,f3,f4,f5);
	dff r30 (e0,clk,rst,y0);
	dff r31 (e1,clk,rst,y1);
	dff r32 (f2,clk,rst,y2);
	dff r33 (f3,clk,rst,y3);
	dff r34 (f4,clk,rst,y4);
	dff r35 (f5,clk,rst,y5);
	dff r36 (e6,clk,rst,y6);
	dff r37 (e7,clk,rst,y7);
endmodule 